module hannwin_f256 (
    input hclk,
    input rst_n,

    //data in 
    input [31:0] data_in,
    input        valid_in,
    output       ready_out,

    //data out
    output [31:0] data_out,
    output        valid_out,
    output        last,         //indicat one frame over, 256 points per frame
    input         ready_in
);

localparam N = 256;
integer i;

reg [31:0] rom_table [N-1:0];
reg [7:0]  counter_in;
wire [31:0] coe;
//-------------------------------------------------------------------------------//
//                               Get right coe                                   //
//===============================================================================//
wire [7:0] counter_in_next;
always @(posedge hclk or negedge rst_n) begin
    if(~rst_n) begin
        counter_in = 8'h00;
    end else begin
        counter_in = counter_in_next;
    end
end
assign counter_in_next = valid_in&ready_out ? counter_in + 1 : counter_in; 
assign coe = rom_table[counter_in];
//-------------------------------------------------------------------------------//
//                        mul       instantiatio                                 //
//===============================================================================//
wire mul_ready_oa, mul_ready_ob;
wire last_in;
assign ready_out = mul_ready_oa & mul_ready_ob;
assign last_in = counter_in==8'hff & valid_in & ready_out;
mul_float32 u0_mul_float32 (
    .aclk(hclk),                                  // input wire aclk
    .aresetn(rst_n),                            // input wire aresetn

    //input data 
    .s_axis_a_tvalid(valid_in),             // input wire s_axis_a_tvalid
    .s_axis_a_tready(mul_ready_oa),            // output wire s_axis_a_tready
    .s_axis_a_tdata(data_in),              // input wire [31 : 0] s_axis_a_tdata
    .s_axis_a_tlast(last_in),              // input wire s_axis_a_tlast
    //rom table 
    .s_axis_b_tvalid(valid_in),            // input wire s_axis_b_tvalid
    .s_axis_b_tready(mul_ready_ob),                      // output wire s_axis_b_tready
    .s_axis_b_tdata(coe),              // input wire [31 : 0] s_axis_b_tdata
    .s_axis_b_tlast(1'b1),              // input wire s_axis_b_tlast

    .m_axis_result_tvalid(valid_out),  // output wire m_axis_result_tvalid
    .m_axis_result_tready(ready_in),  // input wire m_axis_result_tready
    .m_axis_result_tdata(data_out),    // output wire [31 : 0] m_axis_result_tdata
    .m_axis_result_tlast(last)    // output wire m_axis_result_tlast
);


//-------------------------------------------------------------------------------//
//                        initial rom table                                      //
//===============================================================================//
initial begin
    rom_table[0] = 32'b00000000000000000000000000000000;
    rom_table[1] = 32'b00111001000111011110100000000000;
    rom_table[2] = 32'b00111010000111011110001000000000;
    rom_table[3] = 32'b00111010101100011001001100000000;
    rom_table[4] = 32'b00111011000111011100100110000000;
    rom_table[5] = 32'b00111011011101100110111000000000;
    rom_table[6] = 32'b00111011101100010101010100000000;
    rom_table[7] = 32'b00111011111100010011011000000000;
    rom_table[8] = 32'b00111100000111010110100001000000;
    rom_table[9] = 32'b00111100010001110000110001100000;
    rom_table[10] = 32'b00111100011101011000000100000000;
    rom_table[11] = 32'b00111100100101000101111110010000;
    rom_table[12] = 32'b00111100101100000101111101010000;
    rom_table[13] = 32'b00111100110011101011101110010000;
    rom_table[14] = 32'b00111100111011110110111110000000;
    rom_table[15] = 32'b00111101000010010011101100010000;
    rom_table[16] = 32'b00111101000110111110010100010000;
    rom_table[17] = 32'b00111101001011111011001011010000;
    rom_table[18] = 32'b00111101010001001010000101000000;
    rom_table[19] = 32'b00111101010110101010110100111000;
    rom_table[20] = 32'b00111101011100011101001101001000;
    rom_table[21] = 32'b00111101100001010000011111101100;
    rom_table[22] = 32'b00111101100100011010111110011000;
    rom_table[23] = 32'b00111101100111101101111010110100;
    rom_table[24] = 32'b00111101101011001001001100111100;
    rom_table[25] = 32'b00111101101110101100101100001100;
    rom_table[26] = 32'b00111101110010011000001111111000;
    rom_table[27] = 32'b00111101110110001011101110111000;
    rom_table[28] = 32'b00111101111010000110111111110100;
    rom_table[29] = 32'b00111101111110001001111001000000;
    rom_table[30] = 32'b00111110000001001010001000001110;
    rom_table[31] = 32'b00111110000011010010111101111100;
    rom_table[32] = 32'b00111110000101011111011000011010;
    rom_table[33] = 32'b00111110000111101111010010001100;
    rom_table[34] = 32'b00111110001010000010100101101110;
    rom_table[35] = 32'b00111110001100011001001101010110;
    rom_table[36] = 32'b00111110001110110011000011001110;
    rom_table[37] = 32'b00111110010001010000000001011110;
    rom_table[38] = 32'b00111110010011110000000010000000;
    rom_table[39] = 32'b00111110010110010010111110101100;
    rom_table[40] = 32'b00111110011000111000110001001110;
    rom_table[41] = 32'b00111110011011100001010011001010;
    rom_table[42] = 32'b00111110011110001100011110001000;
    rom_table[43] = 32'b00111110100000011101000101101100;
    rom_table[44] = 32'b00111110100001110101001010001100;
    rom_table[45] = 32'b00111110100011001110011001000110;
    rom_table[46] = 32'b00111110100100101000101111000000;
    rom_table[47] = 32'b00111110100110000100001000011100;
    rom_table[48] = 32'b00111110100111100000100001110110;
    rom_table[49] = 32'b00111110101000111101110111101100;
    rom_table[50] = 32'b00111110101010011100000110010110;
    rom_table[51] = 32'b00111110101011111011001010001111;
    rom_table[52] = 32'b00111110101101011010111111101000;
    rom_table[53] = 32'b00111110101110111011100010110110;
    rom_table[54] = 32'b00111110110000011100110000001110;
    rom_table[55] = 32'b00111110110001111110100011111100;
    rom_table[56] = 32'b00111110110011100000111010010001;
    rom_table[57] = 32'b00111110110101000011101111011000;
    rom_table[58] = 32'b00111110110110100110111111011111;
    rom_table[59] = 32'b00111110111000001010100110110010;
    rom_table[60] = 32'b00111110111001101110100001011001;
    rom_table[61] = 32'b00111110111011010010101011100001;
    rom_table[62] = 32'b00111110111100110111000001001101;
    rom_table[63] = 32'b00111110111110011011011110101100;
    rom_table[64] = 32'b00111111000000000000000000000000;
    rom_table[65] = 32'b00111111000000110010010000101011;
    rom_table[66] = 32'b00111111000001100100011111011010;
    rom_table[67] = 32'b00111111000010010110101010010000;
    rom_table[68] = 32'b00111111000011001000101111010100;
    rom_table[69] = 32'b00111111000011111010101100100111;
    rom_table[70] = 32'b00111111000100101100100000010001;
    rom_table[71] = 32'b00111111000101011110001000010101;
    rom_table[72] = 32'b00111111000110001111100010111000;
    rom_table[73] = 32'b00111111000111000000101110000011;
    rom_table[74] = 32'b00111111000111110001100111111010;
    rom_table[75] = 32'b00111111001000100010001110100110;
    rom_table[76] = 32'b00111111001001010010100000001101;
    rom_table[77] = 32'b00111111001010000010011010111001;
    rom_table[78] = 32'b00111111001010110001111100110110;
    rom_table[79] = 32'b00111111001011100001000100001010;
    rom_table[80] = 32'b00111111001100001111101111000110;
    rom_table[81] = 32'b00111111001100111101111011110011;
    rom_table[82] = 32'b00111111001101101011101000100000;
    rom_table[83] = 32'b00111111001110011000110011011110;
    rom_table[84] = 32'b00111111001111000101011010111011;
    rom_table[85] = 32'b00111111001111110001011101001010;
    rom_table[86] = 32'b00111111010000011100111000011110;
    rom_table[87] = 32'b00111111010001000111101011001110;
    rom_table[88] = 32'b00111111010001110001110011101110;
    rom_table[89] = 32'b00111111010010011011010000010101;
    rom_table[90] = 32'b00111111010011000011111111100000;
    rom_table[91] = 32'b00111111010011101011111111101010;
    rom_table[92] = 32'b00111111010100010011001111001100;
    rom_table[93] = 32'b00111111010100111001101100101011;
    rom_table[94] = 32'b00111111010101011111010110100110;
    rom_table[95] = 32'b00111111010110000100001011011110;
    rom_table[96] = 32'b00111111010110101000001001111010;
    rom_table[97] = 32'b00111111010111001011010000100010;
    rom_table[98] = 32'b00111111010111101101011101111110;
    rom_table[99] = 32'b00111111011000001110110000111000;
    rom_table[100] = 32'b00111111011000101111001000000010;
    rom_table[101] = 32'b00111111011001001110100010001010;
    rom_table[102] = 32'b00111111011001101100111110000010;
    rom_table[103] = 32'b00111111011010001010011010011110;
    rom_table[104] = 32'b00111111011010100110110110011001;
    rom_table[105] = 32'b00111111011011000010010000101010;
    rom_table[106] = 32'b00111111011011011100101000001101;
    rom_table[107] = 32'b00111111011011110101111100000011;
    rom_table[108] = 32'b00111111011100001110001011001100;
    rom_table[109] = 32'b00111111011100100101010100101100;
    rom_table[110] = 32'b00111111011100111011010111101100;
    rom_table[111] = 32'b00111111011101010000010011010100;
    rom_table[112] = 32'b00111111011101100100000110110000;
    rom_table[113] = 32'b00111111011101110110110001001111;
    rom_table[114] = 32'b00111111011110001000010010000100;
    rom_table[115] = 32'b00111111011110011000101000100100;
    rom_table[116] = 32'b00111111011110100111110100000110;
    rom_table[117] = 32'b00111111011110110101110100000100;
    rom_table[118] = 32'b00111111011111000010100111111100;
    rom_table[119] = 32'b00111111011111001110001111001111;
    rom_table[120] = 32'b00111111011111011000101001100000;
    rom_table[121] = 32'b00111111011111100001110110010100;
    rom_table[122] = 32'b00111111011111101001110101010110;
    rom_table[123] = 32'b00111111011111110000100110010010;
    rom_table[124] = 32'b00111111011111110110001000110110;
    rom_table[125] = 32'b00111111011111111010011100110111;
    rom_table[126] = 32'b00111111011111111101100010001000;
    rom_table[127] = 32'b00111111011111111111011000100010;
    rom_table[128] = 32'b00111111100000000000000000000000;
    rom_table[129] = 32'b00111111011111111111011000100010;
    rom_table[130] = 32'b00111111011111111101100010001000;
    rom_table[131] = 32'b00111111011111111010011100110110;
    rom_table[132] = 32'b00111111011111110110001000110110;
    rom_table[133] = 32'b00111111011111110000100110010010;
    rom_table[134] = 32'b00111111011111101001110101010110;
    rom_table[135] = 32'b00111111011111100001110110010100;
    rom_table[136] = 32'b00111111011111011000101001011111;
    rom_table[137] = 32'b00111111011111001110001111001110;
    rom_table[138] = 32'b00111111011111000010100111111100;
    rom_table[139] = 32'b00111111011110110101110100000100;
    rom_table[140] = 32'b00111111011110100111110100000101;
    rom_table[141] = 32'b00111111011110011000101000100100;
    rom_table[142] = 32'b00111111011110001000010010000100;
    rom_table[143] = 32'b00111111011101110110110001001110;
    rom_table[144] = 32'b00111111011101100100000110101111;
    rom_table[145] = 32'b00111111011101010000010011010011;
    rom_table[146] = 32'b00111111011100111011010111101100;
    rom_table[147] = 32'b00111111011100100101010100101100;
    rom_table[148] = 32'b00111111011100001110001011001100;
    rom_table[149] = 32'b00111111011011110101111100000010;
    rom_table[150] = 32'b00111111011011011100101000001100;
    rom_table[151] = 32'b00111111011011000010010000101010;
    rom_table[152] = 32'b00111111011010100110110110011000;
    rom_table[153] = 32'b00111111011010001010011010011110;
    rom_table[154] = 32'b00111111011001101100111110000001;
    rom_table[155] = 32'b00111111011001001110100010001001;
    rom_table[156] = 32'b00111111011000101111001000000001;
    rom_table[157] = 32'b00111111011000001110110000110111;
    rom_table[158] = 32'b00111111010111101101011101111100;
    rom_table[159] = 32'b00111111010111001011010000100000;
    rom_table[160] = 32'b00111111010110101000001001111000;
    rom_table[161] = 32'b00111111010110000100001011011110;
    rom_table[162] = 32'b00111111010101011111010110100100;
    rom_table[163] = 32'b00111111010100111001101100101100;
    rom_table[164] = 32'b00111111010100010011001111001101;
    rom_table[165] = 32'b00111111010011101011111111101000;
    rom_table[166] = 32'b00111111010011000011111111011111;
    rom_table[167] = 32'b00111111010010011011010000010100;
    rom_table[168] = 32'b00111111010001110001110011101011;
    rom_table[169] = 32'b00111111010001000111101011001011;
    rom_table[170] = 32'b00111111010000011100111000011111;
    rom_table[171] = 32'b00111111001111110001011101001010;
    rom_table[172] = 32'b00111111001111000101011010111010;
    rom_table[173] = 32'b00111111001110011000110011011100;
    rom_table[174] = 32'b00111111001101101011101000011111;
    rom_table[175] = 32'b00111111001100111101111011110000;
    rom_table[176] = 32'b00111111001100001111101111000011;
    rom_table[177] = 32'b00111111001011100001000100001011;
    rom_table[178] = 32'b00111111001010110001111100110101;
    rom_table[179] = 32'b00111111001010000010011010111001;
    rom_table[180] = 32'b00111111001001010010100000001011;
    rom_table[181] = 32'b00111111001000100010001110100011;
    rom_table[182] = 32'b00111111000111110001100111110111;
    rom_table[183] = 32'b00111111000111000000101110000000;
    rom_table[184] = 32'b00111111000110001111100010111001;
    rom_table[185] = 32'b00111111000101011110001000010100;
    rom_table[186] = 32'b00111111000100101100100000010000;
    rom_table[187] = 32'b00111111000011111010101100100110;
    rom_table[188] = 32'b00111111000011001000101111010010;
    rom_table[189] = 32'b00111111000010010110101010001110;
    rom_table[190] = 32'b00111111000001100100011111010111;
    rom_table[191] = 32'b00111111000000110010010000101011;
    rom_table[192] = 32'b00111111000000000000000000000000;
    rom_table[193] = 32'b00111110111110011011011110101001;
    rom_table[194] = 32'b00111110111100110111000001001010;
    rom_table[195] = 32'b00111110111011010010101011011100;
    rom_table[196] = 32'b00111110111001101110100001010100;
    rom_table[197] = 32'b00111110111000001010100110101100;
    rom_table[198] = 32'b00111110110110100110111111100000;
    rom_table[199] = 32'b00111110110101000011101111010111;
    rom_table[200] = 32'b00111110110011100000111010001110;
    rom_table[201] = 32'b00111110110001111110100011111000;
    rom_table[202] = 32'b00111110110000011100110000001001;
    rom_table[203] = 32'b00111110101110111011100010110010;
    rom_table[204] = 32'b00111110101101011010111111100010;
    rom_table[205] = 32'b00111110101011111011001010001110;
    rom_table[206] = 32'b00111110101010011100000110010110;
    rom_table[207] = 32'b00111110101000111101110111101010;
    rom_table[208] = 32'b00111110100111100000100001110010;
    rom_table[209] = 32'b00111110100110000100001000010111;
    rom_table[210] = 32'b00111110100100101000101110111011;
    rom_table[211] = 32'b00111110100011001110011001000000;
    rom_table[212] = 32'b00111110100001110101001010001100;
    rom_table[213] = 32'b00111110100000011101000101101100;
    rom_table[214] = 32'b00111110011110001100011110000100;
    rom_table[215] = 32'b00111110011011100001010011000110;
    rom_table[216] = 32'b00111110011000111000110001000110;
    rom_table[217] = 32'b00111110010110010010111110100010;
    rom_table[218] = 32'b00111110010011110000000010000010;
    rom_table[219] = 32'b00111110010001010000000001011110;
    rom_table[220] = 32'b00111110001110110011000011001100;
    rom_table[221] = 32'b00111110001100011001001101010010;
    rom_table[222] = 32'b00111110001010000010100101101000;
    rom_table[223] = 32'b00111110000111101111010010000100;
    rom_table[224] = 32'b00111110000101011111011000010010;
    rom_table[225] = 32'b00111110000011010010111101111110;
    rom_table[226] = 32'b00111110000001001010001000001110;
    rom_table[227] = 32'b00111101111110001001111000111100;
    rom_table[228] = 32'b00111101111010000110111111101100;
    rom_table[229] = 32'b00111101110110001011101110110000;
    rom_table[230] = 32'b00111101110010011000001111101100;
    rom_table[231] = 32'b00111101101110101100101100000000;
    rom_table[232] = 32'b00111101101011001001001100111100;
    rom_table[233] = 32'b00111101100111101101111010110100;
    rom_table[234] = 32'b00111101100100011010111110010100;
    rom_table[235] = 32'b00111101100001010000011111100100;
    rom_table[236] = 32'b00111101011100011101001100111000;
    rom_table[237] = 32'b00111101010110101010110100101000;
    rom_table[238] = 32'b00111101010001001010000100110000;
    rom_table[239] = 32'b00111101001011111011001011010000;
    rom_table[240] = 32'b00111101000110111110010100001000;
    rom_table[241] = 32'b00111101000010010011101100010000;
    rom_table[242] = 32'b00111100111011110110111101110000;
    rom_table[243] = 32'b00111100110011101011101101110000;
    rom_table[244] = 32'b00111100101100000101111101000000;
    rom_table[245] = 32'b00111100100101000101111101110000;
    rom_table[246] = 32'b00111100011101011000000100000000;
    rom_table[247] = 32'b00111100010001110000110001100000;
    rom_table[248] = 32'b00111100000111010110100000100000;
    rom_table[249] = 32'b00111011111100010011011000000000;
    rom_table[250] = 32'b00111011101100010101010011000000;
    rom_table[251] = 32'b00111011011101100110111000000000;
    rom_table[252] = 32'b00111011000111011100100100000000;
    rom_table[253] = 32'b00111010101100011001001100000000;
    rom_table[254] = 32'b00111010000111011110001000000000;
    rom_table[255] = 32'b00111001000111011110100000000000;
end






    
endmodule